// *********************************************************************************
// Project Name : CK_riscv
// Author       : Core_kingdom
// Website      : https://blog.csdn.net/weixin_40377195
// Create Time  : 2022-03-12
// File Name    : mux2.v
// Module Name  : mux2
// Called By    :
// Abstract     :
//
// 
// *********************************************************************************
// Modification History:
// Date         By              Version                 Change Description
// -----------------------------------------------------------------------
// 2022-03-12    Macro           1.0                     Original
//  
// *********************************************************************************

module mux2(
    input           sel         ,
    input   [31:0]  data0_in    ,
    input   [31:0]  data1_in    ,

    output  [31:0]  data_out    
);

//=================================================================================
// Parameter declaration
//=================================================================================





//=================================================================================
// Signal declaration
//=================================================================================




//=================================================================================
// Body
//=================================================================================

assign  data_out = (sel == 1'b1) ? data1_in : data0_in;  

endmodule
