// *********************************************************************************
// Project Name : CK_riscv
// Author       : Core_kingdom
// Website      : https://blog.csdn.net/weixin_40377195
// Create Time  : 2022-05-25
// File Name    : CHIP_TOP.v
// Module Name  : CHIP_TOP
// Called By    :
// Abstract     :
//
// 
// *********************************************************************************
// Modification History:
// Date         By              Version                 Change Description
// -----------------------------------------------------------------------
// 2022-05-25    Macro           1.0                     Original
//  
// *********************************************************************************



module CHIP_TOP(
    
    input       sys_clk             ,
    input       sys_rst_n           ,

    output      led_test            

);
//=================================================================================
// Parameter declaration
//=================================================================================


//=================================================================================
// Signal declaration
//=================================================================================


//=================================================================================
// Body
//=================================================================================

riscv_core      u_riscv_core(
    //system signal
    .sys_clk        ( sys_clk       ),
    .sys_rst_n      ( sys_rst_n     ),
    .led_test       ( led_test      )
);

endmodule
